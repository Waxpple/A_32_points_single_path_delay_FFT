module Rom16(
    input clk,
    input rst_n,
    input [5:0] address,
    output reg [21:0] data_real_out,
    output reg [21:0] data_imag_out
);
always@(*)begin
    case (address)
//32 
    6'b100000:begin
//1 
        data_real_out=22'b0000000000000001000000;
//0 
        data_imag_out=22'b0000000000000000000000;
    end
//33 
    6'b100001:begin
//0.98438 
        data_real_out=22'b0000000000000000111111;
//-0.1875 
        data_imag_out=22'b1111111111111111110100;
    end
//34 
    6'b100010:begin
//0.92188 
        data_real_out=22'b0000000000000000111011;
//-0.375 
        data_imag_out=22'b1111111111111111101000;
    end
//35 
    6'b100011:begin
//0.82812 
        data_real_out=22'b0000000000000000110101;
//-0.5625 
        data_imag_out=22'b1111111111111111011100;
    end
//36 
    6'b100100:begin
//0.70312 
        data_real_out=22'b0000000000000000101101;
//-0.70312 
        data_imag_out=22'b1111111111111111010011;
    end
//37 
    6'b100101:begin
//0.5625 
        data_real_out=22'b0000000000000000100100;
//-0.82812 
        data_imag_out=22'b1111111111111111001011;
    end
//38 
    6'b100110:begin
//0.375 
        data_real_out=22'b0000000000000000011000;
//-0.92188 
        data_imag_out=22'b1111111111111111000101;
    end
//39 
    6'b100111:begin
//0.1875 
        data_real_out=22'b0000000000000000001100;
//-0.98438 
        data_imag_out=22'b1111111111111111000001;
    end
//40 
    6'b101000:begin
//0 
        data_real_out=22'b0000000000000000000000;
//-1 
        data_imag_out=22'b1111111111111111000000;
    end
//41 
    6'b101001:begin
//-0.1875 
        data_real_out=22'b1111111111111111110100;
//-0.98438 
        data_imag_out=22'b1111111111111111000001;
    end
//42 
    6'b101010:begin
//-0.375 
        data_real_out=22'b1111111111111111101000;
//-0.92188 
        data_imag_out=22'b1111111111111111000101;
    end
//43 
    6'b101011:begin
//-0.5625 
        data_real_out=22'b1111111111111111011100;
//-0.82812 
        data_imag_out=22'b1111111111111111001011;
    end
//44 
    6'b101100:begin
//-0.70312 
        data_real_out=22'b1111111111111111010011;
//-0.70312 
        data_imag_out=22'b1111111111111111010011;
    end
//45 
    6'b101101:begin
//-0.82812 
        data_real_out=22'b1111111111111111001011;
//-0.5625 
        data_imag_out=22'b1111111111111111011100;
    end
//46 
    6'b101110:begin
//-0.92188 
        data_real_out=22'b1111111111111111000101;
//-0.375 
        data_imag_out=22'b1111111111111111101000;
    end
//47 
    6'b101111:begin
//-0.98438 
        data_real_out=22'b1111111111111111000001;
//-0.1875 
        data_imag_out=22'b1111111111111111110100;
    end
//1 
    default:begin
        data_real_out=23'b0000000000000001000000;
//1 
        data_imag_out=23'b0000000000000000000000;
    end
    endcase
end
endmodule
